Basic RC circuit
r1 1 2 2.0
r2 2 3 3.0
r3 3 0 4.0
r4 3 4 5.0
r5 4 0 6.0
r6 4 0 7.0
*l 1 2 1.0
c 2 0 1.0
vin 1 0  pulse (0 1) ac 1
*.tran  0.1 7.0
.ac dec 10 .01 10
*.plot tran  v(2) i(vin)
.plot ac  vdb(2) xlog
.end
