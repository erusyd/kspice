Basic RC circuit
r 1 2 2.0
c 2 0 1.0
VS 1 0  PWL(15.9N 0.0 16.1n 5.0 31.9n 5.0 32.1n 0.0)
.tran  0.1ns 47ns
.end
